module adjust

fn main() {
	println('Hello World!')
}
