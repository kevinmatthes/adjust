//////////////////////// GNU General Public License 3.0 ////////////////////////
//                                                                            //
// Copyright (C) 2023 Kevin Matthes                                           //
//                                                                            //
// This program is free software: you can redistribute it and/or modify       //
// it under the terms of the GNU General Public License as published by       //
// the Free Software Foundation, either version 3 of the License, or          //
// (at your option) any later version.                                        //
//                                                                            //
// This program is distributed in the hope that it will be useful,            //
// but WITHOUT ANY WARRANTY; without even the implied warranty of             //
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the              //
// GNU General Public License for more details.                               //
//                                                                            //
// You should have received a copy of the GNU General Public License          //
// along with this program.  If not, see <https://www.gnu.org/licenses/>.     //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

module main

import os
import term.ui as terminal

fn main() {
	if os.args.len > 1 {
		if os.args.any(it in ['-h', '--help']) {
			println(help_message)
		} else {
			mut adjust := &Adjust{
				files_to_edit: os.args[1..]
			}

			adjust.window = terminal.init(
				capture_events: true
				event_fn: event_loop
				frame_fn: render
				user_data: adjust
			)

			adjust.window.run()!
		}
	} else {
		println(help_message)
	}
}

////////////////////////////////////////////////////////////////////////////////
